LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY MINUTE IS
	PORT(CLK2, EN2: IN STD_LOGIC;
		 QC: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 CO2: OUT STD_LOGIC;
		 QD: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END MINUTE;

ARCHITECTURE BB OF MINUTE IS
	SIGNAL COUT2, COUT1: STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL CC: STD_LOGIC;
BEGIN
	PROCESS(CLK2, EN2)
	BEGIN
		IF EN2 = '1' THEN
			IF (CLK2'EVENT AND CLK2 = '1') THEN
				IF(COUT2 = 5 AND COUT1 = 8) THEN
				CC <= '1';
				COUT1 <= COUT1 + 1;
				ELSIF (COUT2 = 5 AND COUT1 = 9) THEN
					COUT2 <= "0000";
					COUT1 <= "0000";
					CC <= '0';
				ELSIF (COUT1 = 9) THEN
					COUT2 <= COUT2 + 1;
					COUT1 <= "0000";
					CC <= '0';
				ELSE
					COUT2 <= COUT2;
					COUT1 <= COUT1 + 1;
					CC <= '0';
				END IF;
			END IF;
		END IF;
	END PROCESS;
	CO2 <= CC;
	QC <= COUT2;
	QD <= COUT1;
END BB;
