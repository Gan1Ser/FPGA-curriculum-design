LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY OR_2 IS
	PORT(a,b:IN STD_LOGIC;
		c:OUT STD_LOGIC);
END OR_2;

ARCHITECTURE or2_behavior OF OR_2 IS
BEGIN
	c<=a OR b;
END or2_behavior;