LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY AND_2 IS
	PORT(a,b:IN STD_LOGIC;
		c:OUT STD_LOGIC);
END AND_2;

ARCHITECTURE and2_behavior OF AND_2 IS
BEGIN
	c<=a AND b;
END and2_behavior;