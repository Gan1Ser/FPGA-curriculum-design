LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY HOUR IS
PORT(CLK3, EN3: IN STD_LOGIC;
	 QE,QF : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END HOUR;
ARCHITECTURE BHV OF HOUR IS
	SIGNAL COUNT_SHI, COUNT_GE : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL CLK : STD_LOGIC;
BEGIN 
	CLK <= CLK3 OR (NOT EN3);
	PROCESS(CLK)  	BEGIN
		
			IF CLK'EVENT AND CLK = '1'    THEN
			
				IF COUNT_SHI = "0010" AND COUNT_GE = "0011"		THEN COUNT_SHI <= "0000"; COUNT_GE <= "0000";  -- 24�����������
				ELSIF COUNT_GE < "1001"		THEN COUNT_GE <= COUNT_GE + 1;
				ELSE COUNT_GE <= "0000"; COUNT_SHI <= COUNT_SHI + 1;
				END IF;
			END IF;
		
	QF <=  COUNT_GE;  -- �������
	QE <= COUNT_SHI;
	END PROCESS;
END BHV;