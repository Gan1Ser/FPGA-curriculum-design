LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY FENPIN IS
	PORT(CLK6: IN STD_LOGIC;
		 Q1000: OUT STD_LOGIC;
		 Q1: OUT STD_LOGIC);
END FENPIN;

-- Timer: 16384Hz

ARCHITECTURE CCC_ARC OF FENPIN IS
	SIGNAL X: STD_LOGIC;
BEGIN
	PROCESS(CLK6)
		VARIABLE CNT: INTEGER RANGE 0 TO 32;
	BEGIN
		IF CLK6'EVENT AND CLK6 = '1' THEN
			IF CNT < 31 THEN
				CNT := CNT + 1;
			ELSE
				CNT := 0;
				X <= NOT X;
			END IF;
		END IF;
	END PROCESS;
	
	Q1000 <= X;
	
	PROCESS(X)
		VARIABLE CNT2: INTEGER RANGE 0 TO 256;
		VARIABLE Y: STD_LOGIC;
	BEGIN
		IF X'EVENT AND X = '1' THEN
			IF CNT2 < 255 THEN
				CNT2 := CNT2 + 1;
				Q1 <= '0';
			ELSE
				CNT2 := 0;
				Q1 <= '1';
			END IF;
		END IF;
	END PROCESS;
END CCC_ARC;