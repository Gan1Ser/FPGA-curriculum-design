LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY BEEL_E_CLOCK_VHDL IS 
	PORT(CLK:  IN  STD_LOGIC;
		 SA:   IN  STD_LOGIC;
		 SB:   IN  STD_LOGIC;
		 SC:   IN  STD_LOGIC;
		 INTERRUPT: IN  STD_LOGIC;
		 qw:   OUT STD_LOGIC;
		  r:   OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
	   qout:   OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END BEEL_E_CLOCK_VHDL;

ARCHITECTURE BHV OF  BEEL_E_CLOCK_VHDL IS
	COMPONENT FENPIN 
		PORT(CLK6:  IN  STD_LOGIC;
			Q1000: OUT STD_LOGIC;
			Q1:    OUT STD_LOGIC);
		END COMPONENT;
	
	COMPONENT SECOND IS 
	     PORT(CLK1,EN1:   IN  STD_LOGIC;
	          QA:         OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	          CO1:		  OUT STD_LOGIC;
	          QB:		  OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
	     END COMPONENT;
	COMPONENT MINUTE IS
	     PORT(CLK2,EN2:   IN  STD_LOGIC;
	          QC:         OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	          CO2:		  OUT STD_LOGIC;
	          QD: 		  OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
	     END COMPONENT;
	COMPONENT SelNumber IS 
	     PORT(n1,n2,n3,n4,n5,n6:  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
							  a:  IN  STD_LOGIC_VECTOR(2 DOWNTO 0);    
							qqq:  OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
	     
	     END COMPONENT;
	COMPONENT SelTube   IS
		PORT(M:   IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
			 B:   OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
		END COMPONENT;
	
	COMPONENT HOUR IS
		PORT(CLK3,EN3:   IN  STD_LOGIC;
	          QE:         OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	          QF: 		  OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
	    END COMPONENT;
	
	COMPONENT CNT6 IS
		PORT(CLK5 :IN STD_LOGIC;
	     N:    OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
		END COMPONENT;
		
	COMPONENT OR_2 IS
		PORT(a:   IN STD_LOGIC;
		     b:   IN STD_LOGIC;
		     c:    OUT STD_LOGIC);
		END COMPONENT;
	COMPONENT AND_2 IS 
	    PORT(a:   IN STD_LOGIC;
		     b:   IN STD_LOGIC;
		     c:    OUT STD_LOGIC); 
		END COMPONENT;
		
	COMPONENT DECODER IS
		PORT(a: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		     hex: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
		END COMPONENT;
	
	COMPONENT bell IS
		PORT( CLK4: IN STD_LOGIC;
			  H_SHI, H_GE, M_SHI,M_GE,S_SHI,S_GE:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			  ALARM_OFF: IN STD_LOGIC;
	          speaker:OUT STD_LOGIC);
        END COMPONENT;
     
    SIGNAL m,n,c,h,i,j,z:  STD_LOGIC;
    SIGNAL k,l,e,f,u,v,t:  STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL s:			   STD_LOGIC_VECTOR(2 DOWNTO 0);
    
BEGIN 
	U1:FENPIN  		PORT MAP (CLK6=>CLK,Q1=>h,Q1000=>z);
	U2:SECOND  		PORT MAP (CLK1=>h,EN1=>SC,QA=>k,QB=>l,CO1=>i);
	U3:MINUTE 	    PORT MAP (CLK2=>h,EN2=>m,QC=>e,QD=>f,CO2=>j);
	U4:HOUR    		PORT MAP (CLK3=>h,EN3=>c,QE=>u,QF=>v);
	U5:bell    		PORT MAP (ALARM_OFF=>INTERRUPT,CLK4=>h,H_SHI=>u,H_GE=>v, M_SHI=>e,M_GE=>f,S_SHI=>k,S_GE=>l,speaker=>qw);
    U6:SelNumber	PORT MAP (n1=>u,n2=>v,n3=>e,n4=>f,n5=>k,n6=>l,a=>s,qqq=>t);
    U7:SelTube		PORT MAP (M=>s,B=>r);
    U8:CNT6 		PORT MAP (CLK5=>z,N=>s);
    U9:DECODER		PORT MAP (a=>t,hex=>qout);
    U10:OR_2		PORT MAP (a=>i,b=>SB,c=>m);
    U11:AND_2		PORT MAP (a=>i,b=>j,c=>n);
    U12:OR_2		PORT MAP (a=>n,b=>SA,c=>c);	
     
END BHV;